

module tb;





endmodule;